`timescale 1ns / 1ps



module rep_iter_sel_test;

	// Instantiate the Unit Under Test (UUT)
	rep_iter_selection uut (
	);

	initial begin
		// Initialize Inputs

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here

	end
      
endmodule

