`timescale 1ns / 1ps



module test_repitersel;

	// Instantiate the Unit Under Test (UUT)
	rep_iter_selection uut (
	);

	initial begin
		// Initialize Inputs

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here

	end
      
endmodule

